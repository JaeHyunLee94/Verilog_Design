//full adder using carno map

module full_adder_carno(c1,x,y);

input [3:0] x,y;
output [4:0] c1;
assign c1=x+y;

endmodule


